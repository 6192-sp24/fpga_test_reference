`define TRACE_PORTAL 
`define ConnectalVersion 22.05.23b
`define NumberOfMasters 1
`define PinType Empty
`define PinTypeInclude Misc
`define NumberOfUserTiles 1
`define SlaveDataBusWidth 32
`define SlaveControlAddrWidth 5
`define BurstLenSize 10
`define project_dir $(DTOP)
`define MainClockPeriod 4
`define DerivedClockPeriod 4.000000
`define PcieClockPeriod 4
`define XILINX 1
`define VirtexUltrascale 
`define XilinxUltrascale 
`define PCIE 
`define PCIE3 
`define PcieHostInterface 
`define PhysAddrWidth 40
`define NUMBER_OF_LEDS 2
`define PcieLanes 8
`define CONNECTAL_BITS_DEPENDENCES hw/mkTop.bit
`define CONNECTAL_RUN_SCRIPT $(CONNECTALDIR)/scripts/run.pcietest
`define BOARD_vcu108 
